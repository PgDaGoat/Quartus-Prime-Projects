-- cristinel ababei; 
-- design entity: digital clock, prototyped on Terasic's DE1SoC FPGA board; 
-- EECE-4740 Advanced VHDL Design and FPGAs;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity digital_clock_de1soc is
  Port ( 
    clk_50MHz_external : in STD_LOGIC; -- from crystal quartz oscillator on board; 
    btn_set_seconds: in STD_LOGIC; -- KEY0
    btn_set_minutes : in STD_LOGIC; -- KEY1
    btn_set_hour : in STD_LOGIC; -- KEY2   
    btn_setup_mode : in STD_LOGIC; -- KEY3; keep pressed to setup hour or minutes;
    slide_sw_RESET : in STD_LOGIC; -- reset, SW(0);
    LED_reset : out STD_LOGIC;
    LED_setup_mode : out STD_LOGIC; 
    seven_seg_hour1 : out STD_LOGIC_vector(6 downto 0);
    seven_seg_hour0 : out STD_LOGIC_vector(6 downto 0);
    seven_seg_minutes1 : out STD_LOGIC_vector(6 downto 0);
    seven_seg_minutes0 : out STD_LOGIC_vector(6 downto 0);
    seven_seg_seconds1 : out STD_LOGIC_vector(6 downto 0);
    seven_seg_seconds0 : out STD_LOGIC_vector(6 downto 0)
  );
end digital_clock_de1soc;


architecture my_structural of digital_clock_de1soc is

  COMPONENT clock_counter 
    PORT (
      clk: in std_logic; -- 2MHz main clock;
      reset: in std_logic;
      setup_mode: in std_logic;
      set_hour: in std_logic;
      set_minutes: in std_logic;
      set_seconds: in std_logic;
      hour, minutes, seconds: out std_logic_vector(5 downto 0);
      hour_change, minutes_change, seconds_change: out std_logic
    );
  END COMPONENT;

  COMPONENT bin2bcd 
    PORT (
      clk: in std_logic;
      reset: in std_logic;
      start: in std_logic;
      bin: in std_logic_vector(5 downto 0);
      ready, done_tick: out std_logic;
      bcd1, bcd0: out std_logic_vector(3 downto 0)
    );
  END COMPONENT;
  
  COMPONENT hex_to_sseg
    PORT (
      hex: in std_logic_vector(3 downto 0);
      sseg: out std_logic_vector(6 downto 0)
     );
  END COMPONENT;

  -- Altera PLL; create it with the MegaWizard!
  COMPONENT my_pll 
	port (
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'; --   reset.reset
		outclk_0 : out std_logic         -- outclk0.clk
	);
  end COMPONENT;

  COMPONENT debounce is
    PORT (
      clk, reset: in std_logic;
      sw: in std_logic;
      db: out std_logic
    );
  END COMPONENT;

  -- clocks generated by PLL out of the external clock signal;
  signal clk_2MHz : std_logic;
  
  -- resets;
  signal reset_global : std_logic;
  signal reset_automatic : std_logic;
  signal reset_manual : std_logic;

  -- user controls;
  signal setup_mode, setup_mode_db : std_logic;
  signal set_seconds, set_seconds_db : std_logic;
  signal set_minutes, set_minutes_db : std_logic;
  signal set_hour, set_hour_db : std_logic;
  
  -- other internal signals; bin2bcd is referred to as b2b;
  signal b2b_hour_ready, b2b_hour_start, b2b_hour_done : std_logic;
  signal b2b_minutes_ready, b2b_minutes_start, b2b_minutes_done : std_logic;
  signal b2b_seconds_ready, b2b_seconds_start, b2b_seconds_done : std_logic;
  
  -- hour_bin is the binary value of the current hour; this will
  -- be converted into two BCD digits (bcd1,bcd0); for example,
  -- 000111 gets converted into 07; also,
  -- 001111 gets converted into 15 for 24h display or 03 for AM/PM display;
  -- Note: currently hour is displayed as a number between 1..12; not 0..23;
  signal hour_bin : std_logic_vector(5 downto 0);
  signal hour_bcd1, hour_bcd0 : std_logic_vector(3 downto 0);
  signal minutes_bin : std_logic_vector(5 downto 0);
  signal minutes_bcd1, minutes_bcd0 : std_logic_vector(3 downto 0);
  signal seconds_bin : std_logic_vector(5 downto 0);
  signal seconds_bcd1, seconds_bcd0 : std_logic_vector(3 downto 0); 
 
begin

  
  -- (1) invert push buttons because KEY# on board generates
  -- a signal 111000111; with 1 when not pressed and 0 when pressed/pushed;
  set_seconds <= not btn_set_seconds; -- KEY0;
  set_minutes <= not btn_set_minutes; -- KEY1
  set_hour <= not btn_set_hour; -- KEY2     
  setup_mode <= not btn_setup_mode; -- KEY3
  
  -- (2) debounce slide switch used for manual reset;
  Inst_debounce_reset: debounce PORT MAP(
    clk => clk_50MHz_external,
    reset => '0',
    sw => slide_sw_RESET,
    db => reset_manual
  ); 
  -- first thing when the system is powered on, I should automatically
  -- reset everything for a few clock cycles;
  reset_automatic <= '0';
  reset_global <= (reset_manual or reset_automatic); 

  -- (3) LEDs
  LED_setup_mode <= setup_mode;
  LED_reset <= reset_global;
   
  -- PLL clock: take external 50MHz and slow it down to 2MHz;
  Inst_1_clock_pll: my_pll PORT MAP(
    refclk   => clk_50MHz_external,
		rst      => '0',
		outclk_0 => clk_2MHz
  ); 
  

  -- (4) main clock counter;
  Inst_clock_counter: clock_counter PORT MAP(  
    clk => clk_2MHz,
    reset => reset_global,
    setup_mode => setup_mode,
    set_hour => set_hour,
    set_minutes => set_minutes,
    set_seconds => set_seconds,
    hour => hour_bin,
    minutes => minutes_bin,
    seconds => seconds_bin,
    hour_change => b2b_hour_start, 
    minutes_change => b2b_minutes_start, 
    seconds_change => b2b_seconds_start
  );
 
  
  -- (5) convert the binary values into BCD, which in this case can simply
  -- be converted into 7-segment driving data by interpreting the BCD
  -- as hexadecimal;
  
  -- converter of the hour value into two BCD digits;
  Inst_bin2bcd_hour: bin2bcd PORT MAP(
    clk => clk_2MHz,
    reset => reset_global,
    start => b2b_hour_start,
    bin => hour_bin, -- input binary value to be converted;
    ready => b2b_hour_ready,
    done_tick => b2b_hour_done, -- conversion done; 
    bcd1 => hour_bcd1,
    bcd0 => hour_bcd0
  );
  -- decode the two BCD hour digits into signals needed to drive the 7 segment LED displays;
  Inst_hex_to_sseg_hour1: hex_to_sseg PORT MAP(
    hex => hour_bcd1,
    sseg => seven_seg_hour1
  );
  Inst_hex_to_sseg_hour0: hex_to_sseg PORT MAP(
    hex => hour_bcd0,
    sseg => seven_seg_hour0
  );  

  -- converter of the minutes value into two BCD digits;
  Inst_bin2bcd_minutes: bin2bcd PORT MAP(
    clk => clk_2MHz,
    reset => reset_global,
    start => b2b_minutes_start,
    bin => minutes_bin, -- input binary value to be converted;
    ready => b2b_minutes_ready,
    done_tick => b2b_minutes_done, -- conversion done; 
    bcd1 => minutes_bcd1,
    bcd0 => minutes_bcd0
  ); 
  -- decode the two BCD minutes digits into signals needed to drive the 7 segment LED displays;
  Inst_hex_to_sseg_minutes1: hex_to_sseg PORT MAP(
    hex => minutes_bcd1,
    sseg => seven_seg_minutes1
  );
  Inst_hex_to_sseg_minutes0: hex_to_sseg PORT MAP(
    hex => minutes_bcd0,
    sseg => seven_seg_minutes0
  );  

  -- converter of the seconds value into two BCD digits;
  Inst_bin2bcd_seconds: bin2bcd PORT MAP(
    clk => clk_2MHz,
    reset => reset_global,
    start => b2b_seconds_start, -- high just one cycle;
    bin => seconds_bin, -- input binary value to be converted;
    ready => b2b_seconds_ready, 
    done_tick => b2b_seconds_done, -- conversion done; 
    bcd1 => seconds_bcd1,
    bcd0 => seconds_bcd0
  ); 
  -- decode the two BCD seconds digits into signals needed to drive the 7 
  -- segment LED displays; the two left-most ones on the board;
  Inst_hex_to_sseg_seconds1: hex_to_sseg PORT MAP(
    hex => seconds_bcd1,
    sseg => seven_seg_seconds1
  );
  Inst_hex_to_sseg_seconds0: hex_to_sseg PORT MAP(
    hex => seconds_bcd0,
    sseg => seven_seg_seconds0
  );
 
end my_structural;
